-- This package provides various types useful in testbenches. This version is
-- for VHDL 93
--
-- This Source Code Form is subject to the terms of the Mozilla Public
-- License, v. 2.0. If a copy of the MPL was not distributed with this file,
-- You can obtain one at http://mozilla.org/MPL/2.0/.
--
-- Copyright (c) 2015, Lars Asplund lars.anders.asplund@gmail.com

package test_types is
  subtype shared_natural is natural;
end package test_types;
